module ring_counter ( input clk, reset, output reg [3:0] q);

always@(posedge clk or posedge reset)
  if (reset) 
      q <= 4'b0001;
  else 
      q <= {q[2:0], q[3]};
endmodule
